module uart_fifo #(
    parameter WIDTH = 8,
    parameter DEPTH = 16,
    parameter ALMOST_FULL = 12
) (
    // Read port
    input wire i_rd_en,
    output reg [WIDTH-1:0] o_rd_data,
    output reg o_rd_valid,

    // Write port
    input wire i_wr_en,
    input wire [WIDTH-1:0] i_wr_data,

    // Status
    output wire o_empty,
    output wire o_full,
    output wire o_almostfull,

    input wire i_clk,
    input wire i_rst
);

    localparam ADDR_WIDTH = $clog2(DEPTH);

    reg [WIDTH-1:0] shift_reg [0:DEPTH-1];
    reg [ADDR_WIDTH:0] count = 0; // Declare count to track data in FIFO

    assign o_empty = (count == 0);
    assign o_full = (count == DEPTH);
    assign o_almostfull = (count >= ALMOST_FULL);

    integer i; // Declare integer variable for the shift loop

    always @(posedge i_clk or posedge i_rst) begin
        if (i_rst) begin
            count <= 0;
            o_rd_valid <= 0;
        end else begin
            o_rd_valid <= 0;

            // Write Operation
            if (i_wr_en && !o_full) begin
                shift_reg[count] <= i_wr_data;
                count <= count + 1;
            end

            // Read Operation
            if (i_rd_en && !o_empty) begin
                o_rd_data <= shift_reg[0];
                // Shift data
                for (i = 0; i < DEPTH - 1; i = i + 1) begin
                    shift_reg[i] <= shift_reg[i + 1];
                end
                count <= count - 1;
                o_rd_valid <= 1;
            end
        end
    end
endmodule
